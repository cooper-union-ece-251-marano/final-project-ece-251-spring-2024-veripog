//////////////////////////////////////////////////////////////////////////////////
// The Cooper Union
// ECE 251 Spring 2024
// Engineer: Jaeho Cho & Malek Haddad
// 
//     Create Date: 2023-02-07
//     Module Name: adder
//     Description: simple behavorial adder
//
// Revision: 1.0
//
//////////////////////////////////////////////////////////////////////////////////
`ifndef ADDER
`define ADDER

`timescale 1ns/100ps

module adder
    #(parameter n = 32)(
    input [n-1:0] a,     // n-bit input a
    input [n-1:0] b,     // n-bit input b
    output [n-1:0] sum,  // n-bit sum of a and b
    output carry_out     // Carry out of the addition

);
    // Adding two n-bit numbers
    assign {carry_out, sum} = a + b;

endmodule

`endif // ADDER